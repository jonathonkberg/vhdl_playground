library ieee;
use ieee.std_logic_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity finalcode is
    port(
        clk1,clk2,clk3, reset: in std_logic;
        packet_input: in std_logic_vector(7 downto 0);
        remin: OUT STD_LOGIC_VECTOR (7 downto 0));
        
    end finalcode;
  



architecture hierchical_design of finalcode is
--- COMPONENT DECLARATIONS ---

component dff is
    port(
        D_initial, D: in std_logic;
        clk : in std_logic; 
        Q, Q_n: out std_logic;
        reset : in std_logic
        );
end component;

component dff_8 is
  port(
        D : in std_logic_vector (7 downto 0);
        clk: in std_logic; 
        Q, Q_n: out std_logic_vector (7 downto 0)
    );
end component;

component two_input_xor is
    port(
        input_1, input_2 : in std_logic;
        xor_out : out std_logic
    );
end component;


--- SIGNALS ---

signal f02, f023, feedback: std_logic ;
signal random_number,initial: std_logic_vector (7 downto 0);
signal random_number_out: std_logic_vector (7 downto 0);
signal row_0, row_1, row_2, row_3, row_4, row_5, row_6, row_7,mult_out : std_logic_vector(14 downto 0);
signal ready_0, ready_1, ready_2, ready_3, ready_4, ready_5, ready_6, ready_7, complete : std_logic;
signal start_xor, complete_fsm, populate_rows, reset_rows: std_logic;
signal int1 : std_logic_vector (14 downto 0):= "000000000000000" ;
signal int2 : std_logic_vector (14 downto 0):= "000000000000000";
signal int3 : std_logic_vector (14 downto 0):= "000000000000000" ;
signal int4 : std_logic_vector (14 downto 0):= "000000000000000";
signal int5 : std_logic_vector (14 downto 0):= "000000000000000" ;
signal int6 : std_logic_vector (14 downto 0):= "000000000000000";
signal int7 : std_logic_vector (14 downto 0):= "000000000000000" ;
signal int8 : std_logic_vector (14 downto 0):= "000000000000000";
signal int9 : std_logic_vector (14 downto 0):= "000000000000000" ;
signal int10 : std_logic_vector (14 downto 0):= "000000000000000";
signal int11 : std_logic_vector (14 downto 0):= "000000000000000" ;
signal int12 : std_logic_vector (14 downto 0):= "000000000000000";
signal int13 : std_logic_vector (14 downto 0):= "000000000000000" ;
signal int14 : std_logic_vector (14 downto 0):= "000000000000000";
signal rst : std_logic := '0';
signal flg1 : std_logic := '0';
signal flg2 : std_logic := '0';
signal flg3 : std_logic := '0';
signal flg4 : std_logic := '0';
signal flg5 : std_logic := '0';
signal flg6 : std_logic := '0';
signal flg7 : std_logic := '0';
signal flg : std_logic := '0';
signal Shift_value1 : integer := 0;
signal Shift_value2 : integer := 0;
signal Shift_value3 : integer := 0;
signal Shift_value4 : integer := 0;
signal Shift_value5 : integer := 0;
signal Shift_value6 : integer := 0;
signal Shift_value7 : integer := 0;
signal remin_index  : std_logic_vector (6 downto 0):= "0000000";


--- ARCHITECTURE CONTENT ---

begin

-- initialization process
process(reset)
  begin
    if reset = '1' then
      initial(7) <= '1' after 2 ps;
      initial(6) <= '0' after 2 ps;
      initial(5) <= '1' after 2 ps;
      initial(4) <= '0' after 2 ps;
      initial(3) <= '1' after 2 ps;
      initial(2) <= '0' after 2 ps;
      initial(1) <= '1' after 2 ps;
      initial(0) <= '0' after 2 ps;
    end if;
  end process;


    dff7 : dff
    port map
    (
        D => feedback,
        Q => random_number(7),
        clk => clk1,
        D_initial => initial(7),
        reset => reset
    );
    dff6 : dff
    port map
    (
        D => random_number(7),
        Q => random_number(6),
        clk => clk1,
        D_initial => initial(6),
        reset => reset
    );
    dff5 : dff
    port map
    (
        D => random_number(6),
        Q => random_number(5),
        clk => clk1,
        D_initial => initial(5),
        reset => reset
    );
    dff4 : dff
    port map
    (
        D => random_number(5),
        Q => random_number(4),
        clk => clk1,
        D_initial => initial(4),
        reset => reset
    );
    dff3 : dff
    port map
    (
        D => random_number(4),
        Q => random_number(3),
        clk => clk1,
        D_initial => initial(3),
        reset => reset
    );
    dff2 : dff
    port map
    (
        D => random_number(3),
        Q => random_number(2),
        clk => clk1,
        D_initial => initial(2),
        reset => reset
    );
    dff1 : dff
    port map
    (
        D => random_number(2),
        Q => random_number(1),
        clk => clk1,
        D_initial => initial(1),
        reset => reset
    );
    dff0 : dff
    port map
    (
        D => random_number(1),
        Q => random_number(0),
        clk => clk1,
        D_initial => initial(0),
        reset => reset
    );
    xor_02 : two_input_xor
    port map
    (
        input_1 => random_number(0),
        input_2 => random_number(2),
        xor_out => f02
    );
    xor_023 : two_input_xor
    port map
    (
        input_1 => random_number(3),
        input_2 => f02,
        xor_out => f023
    );
    xor_0234 : two_input_xor
    port map
    (
        input_1 => random_number(4),
        input_2 => f023,
        xor_out => feedback
    );
    dff_out : dff_8
    port map
      (
        D => random_number,
        clk => clk1,
        Q => random_number_out
      );
 --Restart expansion state machine
  -- Full expansion algorithm occurs in one main clock cycle
  -- Signals are re-initialized at restart of state machine
    process(clk2, complete_fsm) is
        begin
          if (clk2 = '1') then
            populate_rows <= '1';
            reset_rows <= '1';
          else
            if(complete_fsm = '1') then
              populate_rows <= '0';
              reset_rows <= '0';
            end if;
          end if;
        end process;
        

-- Row population processes
  -- Processes only populate if populate_rows = 1
  -- Eight rows are populated concurrently
    process(populate_rows) is
      begin
        if(reset_rows = '1') then
          ready_0 <= '0';
          row_0 <= "000000000000000";
        end if;
        if(populate_rows = '1') then
          if (random_number_out(0) = '1') then
            for i in 0 to 7 loop
              row_0(i) <= packet_input(i);
            end loop;
          end if;
          ready_0 <= '1';
        end if;
      end process;

      process(populate_rows) is
        begin
          if(reset_rows = '1') then
            ready_1 <= '0';
            row_1 <= "000000000000000";
          end if;
          if(populate_rows = '1') then
            if (random_number_out(1) = '1') then
              for i in 0 to 7 loop
                row_1(i+1) <= packet_input(i);
              end loop;
            end if;
            ready_1 <= '1';
          end if;
        end process;

        process(populate_rows) is
          begin
            if(reset_rows = '1') then
              ready_2 <= '0';
              row_2 <= "000000000000000";
            end if;
            if(populate_rows = '1') then
              if (random_number_out(2) = '1') then
                for i in 0 to 7 loop
                  row_2(i+2) <= packet_input(i);
                end loop;
              end if;
              ready_2 <= '1';
            end if;
          end process;

          process(populate_rows) is
            begin
              if(reset_rows = '1') then
                ready_3 <= '0';
                row_3 <= "000000000000000";
              end if;
              if(populate_rows = '1') then
                if (random_number_out(3) = '1') then
                  for i in 0 to 7 loop
                    row_3(i+3) <= packet_input(i);
                  end loop;
                end if;
                ready_3 <= '1';
              end if;
            end process;

            process(populate_rows) is
              begin
                if(reset_rows = '1') then
                  ready_4 <= '0';
                  row_4 <= "000000000000000";
                end if;
                if(populate_rows = '1') then
                  if (random_number_out(4) = '1') then
                    for i in 0 to 7 loop
                      row_4(i+4) <= packet_input(i);
                    end loop;
                  end if;
                  ready_4 <= '1';
                end if;
              end process;

              process(populate_rows) is
                begin
                  if(reset_rows = '1') then
                    ready_5 <= '0';
                    row_5 <= "000000000000000";
                  end if;
                  if(populate_rows = '1') then
                    if (random_number_out(5) = '1') then
                      for i in 0 to 7 loop
                        row_5(i+5) <= packet_input(i);
                      end loop;
                    end if;
                    ready_5 <= '1';
                  end if;
                end process;

                process(populate_rows) is
                  begin
                    if(reset_rows = '1') then
                      ready_6 <= '0';
                      row_6 <= "000000000000000";
                    end if;
                    if(populate_rows = '1') then
                      if (random_number_out(6) = '1') then
                        for i in 0 to 7 loop
                          row_6(i+6) <= packet_input(i);
                        end loop;
                      end if;
                      ready_6 <= '1';
                    end if;
                  end process;

                  process(populate_rows) is
                    begin
                      if(reset_rows = '1') then
                        ready_7 <= '0';
                        row_7 <= "000000000000000";
                      end if;
                      if(populate_rows = '1') then
                        if (random_number_out(7) = '1') then
                          for i in 0 to 7 loop
                            row_7(i+7) <= packet_input(i);
                          end loop;
                        end if;
                        ready_7 <= '1';
                      end if;
                    end process;
 
      
        
-- XOR operation
      process(populate_rows, ready_0, ready_1, ready_2, ready_3, ready_4, ready_5, ready_6, ready_7)
        begin
          if (populate_rows = '1') then
            mult_out <= "000000000000000";
            complete_fsm <= '0';
            complete <= '0';
          end if;
          if (ready_0 = '1' and ready_1 = '1' and ready_2 = '1' and ready_3 = '1' and ready_4 = '1' and ready_5 = '1' and ready_6 = '1' and ready_7 = '1') then
            for i in 0 to 14 loop
              mult_out(i) <= (((((((row_0(i) xor row_1(i)) xor row_2(i)) xor row_3(i)) xor row_4(i)) xor row_5(i)) xor row_6(i)) xor row_7(i));
            end loop;
            complete_fsm <= '1';
            complete <= '1';
          end if;
        end process;


check1: process(mult_out,clk3)
   
    begin
      
      if (clk3'event and clk3='1') then
    for i in 14 downto 8 loop
      if mult_out(i) = '1' then 
        flg1 <= '1' ; 
        Shift_value1 <= 14-i ;
        exit ;
     else null  ;
     end if ; 
  end loop ;
 end if; 
end process ; 

Irp_shift1: process (shift_value1)
variable Irp : std_logic_vector (14 downto 0):= "100011011000000" ;

begin 
  int1 <= "000000000000000" ;

  if flg1='1' then
        for i in 14 downto shift_value1 loop
       
        int1(i-shift_value1) <= irp(i) ;
      
  end loop ;
end if;
end process; 

XOR_irp1 :process (int1) 
      
    begin 
   if flg1='1'  then
   for i in 14 downto 0 loop
   int2(i) <= mult_out(i) xor int1(i);
    
end loop;
end if;
end process; 

check2: process(int2,clk3)
   
    begin
      if (clk3'event and clk3='1') then
    for i in 14 downto 8 loop
      if int2(i) = '1' then 
        flg2 <= '1' ;
        Shift_value2 <= 14-i ;
        exit ;
     else flg2 <= '0' ; 
     end if ; 
  end loop ;
end if;
end process ; 

Irp_shift2: process (Shift_value2)
variable Irp : std_logic_vector (14 downto 0):= "100011011000000" ;

begin 
  int3 <= "000000000000000" ;
  --flg1 <= '0';
  --if (clk'event and clk='1') then
  if flg2='1' then
        for i in 14 downto shift_value2 loop
       
        int3(i-shift_value2) <= irp(i) ;
      
  end loop ;
  
end if;
end process; 

XOR_irp2 :process (int3) 
      
    begin 
  --if (clk'event and clk='1') and  
   if flg2='1' then
   for i in 14 downto 0 loop
   int4(i) <= int2(i) xor int3(i);
    
end loop;
end if;
end process;

check3: process(int4,clk3)
   
    begin
     if (clk3'event and clk3='1') then 
    for i in 14 downto 8 loop
      if int4(i) = '1' then 
        flg3 <= '1' ;
        Shift_value3 <= 14-i ;
        exit ;
     else flg3 <= '0' ; 
     end if ; 
  end loop ;
end if;
end process ; 

Irp_shift3: process (Shift_value3)
variable Irp : std_logic_vector (14 downto 0):= "100011011000000" ;

begin 
  int5 <= "000000000000000" ;
 -- if (clk'event and clk='1') then
    if flg3='1' then
        for i in 14 downto shift_value3 loop
       
        int5(i-shift_value3) <= irp(i) ;
      
  end loop ;
  
end if;
end process; 

XOR_irp3 :process (int5) 
      
    begin 
   --if (clk'event and clk='1') and
    if flg3='1'  then
   for i in 14 downto 0 loop
   int6(i) <= int4(i) xor int5(i);
    
end loop;
end if;
end process; 

check4: process(int6,clk3)
   
    begin
    if (clk3'event and clk3='1') then  
    for i in 14 downto 8 loop
      if int6(i) = '1' then 
        flg4 <= '1' ;
        Shift_value4 <= 14-i ;
        exit ;
     else flg4 <= '0' ;
     end if ; 
  end loop ;
end if;
end process ; 

Irp_shift4: process (Shift_value4)
variable Irp : std_logic_vector (14 downto 0):= "100011011000000" ;

begin 
  int7 <= "000000000000000" ;
  --if (clk'event and clk='1') then
     if flg4='1' then
        for i in 14 downto shift_value4 loop
       
        int7(i-shift_value4) <= irp(i) ;
      
  end loop ;
 
end if;
end process; 

XOR_irp4 :process (int7) 
      
    begin 
   --if (clk'event and clk='1') and 
   if flg4='1'  then
   for i in 14 downto 0 loop
   int8(i) <= int6(i) xor int7(i);
    
end loop;
end if;
end process;

check5: process(int8,clk3)
   
    begin
      if (clk3'event and clk3='1') then
    for i in 14 downto 8 loop
      if int8(i) = '1' then 
        flg5 <= '1' ;
        Shift_value5 <= 14-i ;
        exit ;
     else flg5 <= '0' ; 
     end if ; 
  end loop ;
end if;
end process ; 

Irp_shift5: process (Shift_value5)
variable Irp : std_logic_vector (14 downto 0):= "100011011000000" ;

begin 
  int9 <= "000000000000000" ;
  --if (clk'event and clk='1') then
     if flg5='1' then
        for i in 14 downto shift_value5 loop
       
        int9(i-shift_value5) <= irp(i) ;
      
  end loop ;
 
end if;
end process; 

XOR_irp5 :process (int9) 
      
    begin 
  -- if (clk'event and clk='1') and
   if flg5='1'  then
   for i in 14 downto 0 loop
   int10(i) <= int8(i) xor int9(i);
    
end loop;
end if;
end process;
check6: process(int10,clk3)
   
    begin
     if (clk3'event and clk3='1') then 
    for i in 14 downto 8 loop
      if int10(i) = '1' then 
        flg6 <= '1' ;
        Shift_value6 <= 14-i ;
        exit ;
     else flg6 <= '0' ; 
     end if ; 
  end loop ;
end if;
end process ; 

Irp_shift6: process (Shift_value6)
variable Irp : std_logic_vector (14 downto 0):= "100011011000000" ;

begin 
  int11 <= "000000000000000" ;
  --if (clk'event and clk='1') then
     if flg6='1' then
        for i in 14 downto shift_value6 loop
       
        int11(i-shift_value6) <= irp(i) ;
      
  end loop ;
  
end if;
end process; 

XOR_irp6 :process (int11) 
      
    begin 
   --if (clk'event and clk='1') and
   if flg6='1'  then
   for i in 14 downto 0 loop
   int12(i) <= int10(i) xor int11(i);
    
end loop;
end if;
end process; 


 check7: process(int12,clk3)
   
    begin
     if (clk3'event and clk3='1') then 
    for i in 14 downto 8 loop
      if int12(i) = '1' then 
        flg7 <= '1' ;
        Shift_value7 <= 14-i ;
        exit ;
     else flg7 <= '0' ; 
     end if ; 
  end loop ;
end if;
end process ; 

Irp_shift7: process (Shift_value7)
variable Irp : std_logic_vector (14 downto 0):= "100011011000000" ;

begin 
  int13 <= "000000000000000" ;
  --if (clk'event and clk='1') then
     if flg7='1' then
        for i in 14 downto shift_value7 loop
       
        int13(i-shift_value7) <= irp(i) ;
      
  end loop ;
  
end if;
end process; 

XOR_irp7 :process (int13) 
      
    begin 
   --if (clk'event and clk='1') and 
   if flg7='1'  then
   for i in 14 downto 0 loop
   int14(i) <= int12(i) xor int13(i);
    
end loop;
end if;
end process; 

concat :process (clk3) 
      
    begin 
      remin_index  <=  flg1 & flg2 & flg3 & flg4 & flg5 & flg6 & flg7  ;

end process; 

Reminder :process (remin_index) 
      
    begin 

 case remin_index is
            when "0000000" =>
                remin <= mult_out(7 downto 0); 
            when "1000000" =>
                remin <= int2(7 downto 0);
            when "1100000" =>
                remin <= int4(7 downto 0);
            when "1110000" =>
                remin <= int6(7 downto 0);
            when "1111000" =>
                 remin <= int8(7 downto 0);
            when "1111100" =>
                 remin <= int10(7 downto 0);
            when "1111110" =>
                 remin <= int12(7 downto 0);
            when others => -- 'U', 'X', '-', etc.
                remin <= int14(7 downto 0) ;
        end case;
 

end process; 


 end hierchical_design;

