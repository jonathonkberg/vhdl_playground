//
// Verilog description for cell galois_expand, 
// Thu May  4 21:52:18 2023
//
// LeonardoSpectrum Level 3, 2011a.4 
//


module galois_expand ( clk, packet_input, random_num_input, mult_out, complete
                        ) ;

    input clk ;
    input [7:0]packet_input ;
    input [7:0]random_num_input ;
    output [14:0]mult_out ;
    output complete ;

    wire nx2453, row_0_0, reset_rows, ready_1, nx16, nx24, nx26, row_0_1, nx36, 
         row_1_1, nx44, nx54, row_0_2, nx64, row_1_2, nx72, row_2_2, nx82, nx90, 
         nx92, row_0_3, nx102, row_1_3, nx110, row_2_3, nx120, nx128, row_3_3, 
         nx130, nx140, row_4_4, nx148, row_0_4, nx158, row_1_4, nx166, row_2_4, 
         nx176, row_3_4, nx184, nx196, nx198, row_0_5, nx208, row_1_5, nx216, 
         row_2_5, nx226, row_3_5, nx234, row_4_5, nx246, row_5_5, nx254, nx266, 
         row_0_6, nx276, row_1_6, nx284, row_2_6, nx294, row_3_6, nx302, row_6_6, 
         nx314, row_4_6, nx322, row_5_6, nx330, nx340, nx342, nx344, row_0_7, 
         nx354, row_1_7, nx362, row_2_7, nx372, row_3_7, nx380, row_4_7, nx392, 
         row_5_7, nx400, row_6_7, nx410, row_7_7, nx418, nx432, row_1_8, nx440, 
         row_2_8, nx448, row_3_8, nx458, row_4_8, nx466, row_7_8, nx478, row_5_8, 
         nx486, row_6_8, nx494, nx504, nx506, nx508, row_2_9, nx516, row_3_9, 
         nx524, row_4_9, nx534, row_5_9, nx542, row_6_9, nx554, row_7_9, nx562, 
         nx574, row_7_10, nx582, row_3_10, nx590, row_4_10, nx598, row_5_10, 
         nx608, row_6_10, nx616, nx628, nx630, row_4_11, nx638, row_5_11, nx646, 
         row_6_11, nx656, nx664, row_7_11, nx666, nx676, row_5_12, nx684, 
         row_6_12, nx692, row_7_12, nx702, nx710, nx712, row_6_13, nx720, 
         row_7_13, nx728, nx738, row_7_14, nx746, nx754, nx2506, nx2511, nx2515, 
         nx2524, nx2528, nx2538, nx2541, nx2545, nx2562, nx2564, nx2568, nx2572, 
         nx2580, nx2582, nx2584, nx2588, nx2592, nx2598, nx2609, nx2611, nx2615, 
         nx2619, nx2630, nx2638, nx2640, nx2642, nx2646, nx2650, nx2656, nx2658, 
         nx2664, nx2675, nx2677, nx2683, nx2692, nx2700, nx2702, nx2704, nx2710, 
         nx2716, nx2727, nx2729, nx2735, nx2743, nx2746, nx2759, nx2769, nx2784, 
         nx2786, nx2788, nx2790, nx2792, nx2794, nx2796, nx2798, nx2800, nx2802, 
         nx2804, nx2806, nx2808, nx2810, nx2814, nx2816, nx2818, nx2820, nx2822, 
         nx2826, nx2830, nx2832, nx2836, nx2840, nx2846, nx2848, nx2852, nx2856, 
         nx2860, nx2862, nx2864, nx5, nx2870, nx2872, nx2874, nx2876;



    fake_gnd ix2454 (.Y (nx2453)) ;
    latch lat_mult_out_0 (.Q (mult_out[0]), .D (nx24), .CLK (nx2814)) ;
    latch lat_row_0_0 (.Q (row_0_0), .D (nx16), .CLK (nx2860)) ;
    nand02 ix2507 (.Y (nx2506), .A0 (packet_input[0]), .A1 (nx2860)) ;
    latch lat_mult_out_1 (.Q (mult_out[1]), .D (nx54), .CLK (nx2814)) ;
    xnor2 ix2512 (.Y (nx2511), .A0 (row_0_1), .A1 (row_1_1)) ;
    latch lat_row_0_1 (.Q (row_0_1), .D (nx36), .CLK (nx2786)) ;
    nand02 ix2516 (.Y (nx2515), .A0 (packet_input[1]), .A1 (nx2860)) ;
    latch lat_row_1_1 (.Q (row_1_1), .D (nx44), .CLK (nx2786)) ;
    latch lat_mult_out_2 (.Q (mult_out[2]), .D (nx92), .CLK (nx2814)) ;
    xnor2 ix91 (.Y (nx90), .A0 (nx2524), .A1 (row_2_2)) ;
    xnor2 ix2525 (.Y (nx2524), .A0 (row_0_2), .A1 (row_1_2)) ;
    latch lat_row_0_2 (.Q (row_0_2), .D (nx64), .CLK (nx2786)) ;
    nand02 ix2529 (.Y (nx2528), .A0 (packet_input[2]), .A1 (nx2786)) ;
    latch lat_row_1_2 (.Q (row_1_2), .D (nx72), .CLK (nx2786)) ;
    latch lat_row_2_2 (.Q (row_2_2), .D (nx82), .CLK (nx2786)) ;
    latch lat_mult_out_3 (.Q (mult_out[3]), .D (nx140), .CLK (nx2814)) ;
    xnor2 ix2539 (.Y (nx2538), .A0 (nx128), .A1 (row_3_3)) ;
    xnor2 ix129 (.Y (nx128), .A0 (nx2541), .A1 (row_2_3)) ;
    xnor2 ix2542 (.Y (nx2541), .A0 (row_0_3), .A1 (row_1_3)) ;
    latch lat_row_0_3 (.Q (row_0_3), .D (nx102), .CLK (nx2788)) ;
    nand02 ix2546 (.Y (nx2545), .A0 (packet_input[3]), .A1 (nx2788)) ;
    latch lat_row_1_3 (.Q (row_1_3), .D (nx110), .CLK (nx2788)) ;
    latch lat_row_2_3 (.Q (row_2_3), .D (nx120), .CLK (nx2788)) ;
    latch lat_row_3_3 (.Q (row_3_3), .D (nx130), .CLK (nx2788)) ;
    latch lat_mult_out_4 (.Q (mult_out[4]), .D (nx198), .CLK (nx2814)) ;
    xnor2 ix197 (.Y (nx196), .A0 (row_4_4), .A1 (nx2562)) ;
    latch lat_row_4_4 (.Q (row_4_4), .D (nx148), .CLK (nx2788)) ;
    xnor2 ix2563 (.Y (nx2562), .A0 (nx2564), .A1 (nx2572)) ;
    xnor2 ix2565 (.Y (nx2564), .A0 (row_0_4), .A1 (row_1_4)) ;
    latch lat_row_0_4 (.Q (row_0_4), .D (nx158), .CLK (nx2862)) ;
    nand02 ix2569 (.Y (nx2568), .A0 (packet_input[4]), .A1 (nx2862)) ;
    latch lat_row_1_4 (.Q (row_1_4), .D (nx166), .CLK (nx2862)) ;
    xnor2 ix2573 (.Y (nx2572), .A0 (row_2_4), .A1 (row_3_4)) ;
    latch lat_row_2_4 (.Q (row_2_4), .D (nx176), .CLK (nx2862)) ;
    latch lat_row_3_4 (.Q (row_3_4), .D (nx184), .CLK (nx2862)) ;
    latch lat_mult_out_5 (.Q (mult_out[5]), .D (nx266), .CLK (nx2814)) ;
    xnor2 ix2581 (.Y (nx2580), .A0 (nx2582), .A1 (nx2598)) ;
    xnor2 ix2583 (.Y (nx2582), .A0 (nx2584), .A1 (nx2592)) ;
    xnor2 ix2585 (.Y (nx2584), .A0 (row_0_5), .A1 (row_1_5)) ;
    latch lat_row_0_5 (.Q (row_0_5), .D (nx208), .CLK (nx2792)) ;
    nand02 ix2589 (.Y (nx2588), .A0 (packet_input[5]), .A1 (nx2862)) ;
    latch lat_row_1_5 (.Q (row_1_5), .D (nx216), .CLK (nx2792)) ;
    xnor2 ix2593 (.Y (nx2592), .A0 (row_2_5), .A1 (row_3_5)) ;
    latch lat_row_2_5 (.Q (row_2_5), .D (nx226), .CLK (nx2792)) ;
    latch lat_row_3_5 (.Q (row_3_5), .D (nx234), .CLK (nx2792)) ;
    xnor2 ix2599 (.Y (nx2598), .A0 (row_4_5), .A1 (row_5_5)) ;
    latch lat_row_4_5 (.Q (row_4_5), .D (nx246), .CLK (nx2792)) ;
    latch lat_row_5_5 (.Q (row_5_5), .D (nx254), .CLK (nx2792)) ;
    latch lat_mult_out_6 (.Q (mult_out[6]), .D (nx344), .CLK (nx2816)) ;
    xnor2 ix343 (.Y (nx342), .A0 (nx2609), .A1 (nx340)) ;
    xnor2 ix2610 (.Y (nx2609), .A0 (nx2611), .A1 (nx2619)) ;
    xnor2 ix2612 (.Y (nx2611), .A0 (row_0_6), .A1 (row_1_6)) ;
    latch lat_row_0_6 (.Q (row_0_6), .D (nx276), .CLK (nx2794)) ;
    nand02 ix2616 (.Y (nx2615), .A0 (packet_input[6]), .A1 (nx2794)) ;
    latch lat_row_1_6 (.Q (row_1_6), .D (nx284), .CLK (nx2794)) ;
    xnor2 ix2620 (.Y (nx2619), .A0 (row_2_6), .A1 (row_3_6)) ;
    latch lat_row_2_6 (.Q (row_2_6), .D (nx294), .CLK (nx2794)) ;
    latch lat_row_3_6 (.Q (row_3_6), .D (nx302), .CLK (nx2794)) ;
    xnor2 ix341 (.Y (nx340), .A0 (row_6_6), .A1 (nx2630)) ;
    latch lat_row_6_6 (.Q (row_6_6), .D (nx314), .CLK (nx2794)) ;
    xnor2 ix2631 (.Y (nx2630), .A0 (row_4_6), .A1 (row_5_6)) ;
    latch lat_row_4_6 (.Q (row_4_6), .D (nx322), .CLK (nx2796)) ;
    latch lat_row_5_6 (.Q (row_5_6), .D (nx330), .CLK (nx2796)) ;
    latch lat_mult_out_7 (.Q (mult_out[7]), .D (nx432), .CLK (nx2816)) ;
    xnor2 ix2639 (.Y (nx2638), .A0 (nx2640), .A1 (nx2656)) ;
    xnor2 ix2641 (.Y (nx2640), .A0 (nx2642), .A1 (nx2650)) ;
    xnor2 ix2643 (.Y (nx2642), .A0 (row_0_7), .A1 (row_1_7)) ;
    latch lat_row_0_7 (.Q (row_0_7), .D (nx354), .CLK (nx2796)) ;
    nand02 ix2647 (.Y (nx2646), .A0 (packet_input[7]), .A1 (nx2796)) ;
    latch lat_row_1_7 (.Q (row_1_7), .D (nx362), .CLK (nx2796)) ;
    xnor2 ix2651 (.Y (nx2650), .A0 (row_2_7), .A1 (row_3_7)) ;
    latch lat_row_2_7 (.Q (row_2_7), .D (nx372), .CLK (nx2796)) ;
    latch lat_row_3_7 (.Q (row_3_7), .D (nx380), .CLK (nx2798)) ;
    xnor2 ix2657 (.Y (nx2656), .A0 (nx2658), .A1 (nx2664)) ;
    xnor2 ix2659 (.Y (nx2658), .A0 (row_4_7), .A1 (row_5_7)) ;
    latch lat_row_4_7 (.Q (row_4_7), .D (nx392), .CLK (nx2798)) ;
    latch lat_row_5_7 (.Q (row_5_7), .D (nx400), .CLK (nx2798)) ;
    xnor2 ix2665 (.Y (nx2664), .A0 (row_6_7), .A1 (row_7_7)) ;
    latch lat_row_6_7 (.Q (row_6_7), .D (nx410), .CLK (nx2798)) ;
    latch lat_row_7_7 (.Q (row_7_7), .D (nx418), .CLK (nx2798)) ;
    latch lat_mult_out_8 (.Q (mult_out[8]), .D (nx508), .CLK (nx2816)) ;
    xnor2 ix507 (.Y (nx506), .A0 (nx2675), .A1 (nx504)) ;
    xnor2 ix2676 (.Y (nx2675), .A0 (nx2677), .A1 (nx2683)) ;
    xnor2 ix2678 (.Y (nx2677), .A0 (row_1_8), .A1 (row_2_8)) ;
    latch lat_row_1_8 (.Q (row_1_8), .D (nx440), .CLK (nx2798)) ;
    latch lat_row_2_8 (.Q (row_2_8), .D (nx448), .CLK (nx2800)) ;
    xnor2 ix2684 (.Y (nx2683), .A0 (row_3_8), .A1 (row_4_8)) ;
    latch lat_row_3_8 (.Q (row_3_8), .D (nx458), .CLK (nx2800)) ;
    latch lat_row_4_8 (.Q (row_4_8), .D (nx466), .CLK (nx2800)) ;
    xnor2 ix505 (.Y (nx504), .A0 (row_7_8), .A1 (nx2692)) ;
    latch lat_row_7_8 (.Q (row_7_8), .D (nx478), .CLK (nx2800)) ;
    xnor2 ix2693 (.Y (nx2692), .A0 (row_5_8), .A1 (row_6_8)) ;
    latch lat_row_5_8 (.Q (row_5_8), .D (nx486), .CLK (nx2800)) ;
    latch lat_row_6_8 (.Q (row_6_8), .D (nx494), .CLK (nx2800)) ;
    latch lat_mult_out_9 (.Q (mult_out[9]), .D (nx574), .CLK (nx2816)) ;
    xnor2 ix2701 (.Y (nx2700), .A0 (nx2702), .A1 (nx2716)) ;
    xnor2 ix2703 (.Y (nx2702), .A0 (nx2704), .A1 (nx2710)) ;
    xnor2 ix2705 (.Y (nx2704), .A0 (row_2_9), .A1 (row_3_9)) ;
    latch lat_row_2_9 (.Q (row_2_9), .D (nx516), .CLK (nx2802)) ;
    latch lat_row_3_9 (.Q (row_3_9), .D (nx524), .CLK (nx2802)) ;
    xnor2 ix2711 (.Y (nx2710), .A0 (row_4_9), .A1 (row_5_9)) ;
    latch lat_row_4_9 (.Q (row_4_9), .D (nx534), .CLK (nx2802)) ;
    latch lat_row_5_9 (.Q (row_5_9), .D (nx542), .CLK (nx2802)) ;
    xnor2 ix2717 (.Y (nx2716), .A0 (row_6_9), .A1 (row_7_9)) ;
    latch lat_row_6_9 (.Q (row_6_9), .D (nx554), .CLK (nx2802)) ;
    latch lat_row_7_9 (.Q (row_7_9), .D (nx562), .CLK (nx2802)) ;
    latch lat_mult_out_10 (.Q (mult_out[10]), .D (nx630), .CLK (nx2816)) ;
    xnor2 ix629 (.Y (nx628), .A0 (row_7_10), .A1 (nx2727)) ;
    latch lat_row_7_10 (.Q (row_7_10), .D (nx582), .CLK (nx2804)) ;
    xnor2 ix2728 (.Y (nx2727), .A0 (nx2729), .A1 (nx2735)) ;
    xnor2 ix2730 (.Y (nx2729), .A0 (row_3_10), .A1 (row_4_10)) ;
    latch lat_row_3_10 (.Q (row_3_10), .D (nx590), .CLK (nx2804)) ;
    latch lat_row_4_10 (.Q (row_4_10), .D (nx598), .CLK (nx2804)) ;
    xnor2 ix2736 (.Y (nx2735), .A0 (row_5_10), .A1 (row_6_10)) ;
    latch lat_row_5_10 (.Q (row_5_10), .D (nx608), .CLK (nx2804)) ;
    latch lat_row_6_10 (.Q (row_6_10), .D (nx616), .CLK (nx2804)) ;
    latch lat_mult_out_11 (.Q (mult_out[11]), .D (nx676), .CLK (nx2816)) ;
    xnor2 ix2744 (.Y (nx2743), .A0 (nx664), .A1 (row_7_11)) ;
    xnor2 ix665 (.Y (nx664), .A0 (nx2746), .A1 (row_6_11)) ;
    xnor2 ix2747 (.Y (nx2746), .A0 (row_4_11), .A1 (row_5_11)) ;
    latch lat_row_4_11 (.Q (row_4_11), .D (nx638), .CLK (nx2804)) ;
    latch lat_row_5_11 (.Q (row_5_11), .D (nx646), .CLK (nx2806)) ;
    latch lat_row_6_11 (.Q (row_6_11), .D (nx656), .CLK (nx2806)) ;
    latch lat_row_7_11 (.Q (row_7_11), .D (nx666), .CLK (nx2806)) ;
    latch lat_mult_out_12 (.Q (mult_out[12]), .D (nx712), .CLK (nx26)) ;
    xnor2 ix711 (.Y (nx710), .A0 (nx2759), .A1 (row_7_12)) ;
    xnor2 ix2760 (.Y (nx2759), .A0 (row_5_12), .A1 (row_6_12)) ;
    latch lat_row_5_12 (.Q (row_5_12), .D (nx684), .CLK (nx2806)) ;
    latch lat_row_6_12 (.Q (row_6_12), .D (nx692), .CLK (nx2806)) ;
    latch lat_row_7_12 (.Q (row_7_12), .D (nx702), .CLK (nx2806)) ;
    latch lat_mult_out_13 (.Q (mult_out[13]), .D (nx738), .CLK (nx26)) ;
    xnor2 ix2770 (.Y (nx2769), .A0 (row_6_13), .A1 (row_7_13)) ;
    latch lat_row_6_13 (.Q (row_6_13), .D (nx720), .CLK (nx2808)) ;
    latch lat_row_7_13 (.Q (row_7_13), .D (nx728), .CLK (nx2808)) ;
    latch lat_mult_out_14 (.Q (mult_out[14]), .D (nx754), .CLK (nx26)) ;
    latch lat_row_7_14 (.Q (row_7_14), .D (nx746), .CLK (nx2808)) ;
    inv01 ix2783 (.Y (nx2784), .A (nx2864)) ;
    inv01 ix2785 (.Y (nx2786), .A (nx2864)) ;
    inv01 ix2787 (.Y (nx2788), .A (nx2864)) ;
    inv01 ix2789 (.Y (nx2790), .A (nx2864)) ;
    inv01 ix2791 (.Y (nx2792), .A (nx2864)) ;
    inv01 ix2793 (.Y (nx2794), .A (nx2820)) ;
    inv01 ix2795 (.Y (nx2796), .A (nx2820)) ;
    inv01 ix2797 (.Y (nx2798), .A (nx2820)) ;
    inv01 ix2799 (.Y (nx2800), .A (nx2820)) ;
    inv01 ix2801 (.Y (nx2802), .A (nx2820)) ;
    inv01 ix2803 (.Y (nx2804), .A (nx2820)) ;
    inv01 ix2805 (.Y (nx2806), .A (nx2822)) ;
    inv01 ix2807 (.Y (nx2808), .A (nx2822)) ;
    inv01 ix2809 (.Y (nx2810), .A (nx2876)) ;
    inv01 ix2817 (.Y (nx2818), .A (reset_rows)) ;
    inv01 ix2819 (.Y (nx2820), .A (reset_rows)) ;
    inv01 ix2821 (.Y (nx2822), .A (reset_rows)) ;
    inv01 ix2825 (.Y (nx2826), .A (nx2874)) ;
    nand02 ix2829 (.Y (nx2830), .A0 (packet_input[0]), .A1 (nx2784)) ;
    nand02 ix2831 (.Y (nx2832), .A0 (packet_input[1]), .A1 (nx2784)) ;
    nand02 ix2835 (.Y (nx2836), .A0 (packet_input[2]), .A1 (nx2786)) ;
    nand02 ix2839 (.Y (nx2840), .A0 (packet_input[3]), .A1 (nx2788)) ;
    nand02 ix2845 (.Y (nx2846), .A0 (packet_input[4]), .A1 (nx2790)) ;
    nand02 ix2847 (.Y (nx2848), .A0 (packet_input[5]), .A1 (nx2790)) ;
    nand02 ix2851 (.Y (nx2852), .A0 (packet_input[6]), .A1 (nx2794)) ;
    nand02 ix2855 (.Y (nx2856), .A0 (packet_input[7]), .A1 (nx2796)) ;
    inv01 ix2859 (.Y (nx2860), .A (nx2818)) ;
    inv01 ix2861 (.Y (nx2862), .A (nx2818)) ;
    inv01 ix2863 (.Y (nx2864), .A (reset_rows)) ;
    nor02ii ix25 (.Y (nx24), .A0 (nx2876), .A1 (row_0_0)) ;
    nor02ii ix17 (.Y (nx16), .A0 (nx2830), .A1 (random_num_input[0])) ;
    or02 ix27 (.Y (nx26), .A0 (reset_rows), .A1 (nx2874)) ;
    nor02ii ix55 (.Y (nx54), .A0 (nx2511), .A1 (nx2874)) ;
    nor02ii ix37 (.Y (nx36), .A0 (nx2832), .A1 (random_num_input[0])) ;
    nor02ii ix45 (.Y (nx44), .A0 (nx2830), .A1 (random_num_input[1])) ;
    nor02ii ix93 (.Y (nx92), .A0 (nx2876), .A1 (nx90)) ;
    nor02ii ix65 (.Y (nx64), .A0 (nx2836), .A1 (random_num_input[0])) ;
    nor02ii ix73 (.Y (nx72), .A0 (nx2832), .A1 (random_num_input[1])) ;
    nor02ii ix83 (.Y (nx82), .A0 (nx2830), .A1 (random_num_input[2])) ;
    nor02ii ix141 (.Y (nx140), .A0 (nx2538), .A1 (nx2874)) ;
    nor02ii ix103 (.Y (nx102), .A0 (nx2840), .A1 (random_num_input[0])) ;
    nor02ii ix111 (.Y (nx110), .A0 (nx2836), .A1 (random_num_input[1])) ;
    nor02ii ix121 (.Y (nx120), .A0 (nx2832), .A1 (random_num_input[2])) ;
    nor02ii ix131 (.Y (nx130), .A0 (nx2830), .A1 (random_num_input[3])) ;
    nor02ii ix199 (.Y (nx198), .A0 (nx2876), .A1 (nx196)) ;
    nor02ii ix149 (.Y (nx148), .A0 (nx2830), .A1 (random_num_input[4])) ;
    nor02ii ix159 (.Y (nx158), .A0 (nx2846), .A1 (random_num_input[0])) ;
    nor02ii ix167 (.Y (nx166), .A0 (nx2840), .A1 (random_num_input[1])) ;
    nor02ii ix177 (.Y (nx176), .A0 (nx2836), .A1 (random_num_input[2])) ;
    nor02ii ix185 (.Y (nx184), .A0 (nx2832), .A1 (random_num_input[3])) ;
    nor02ii ix267 (.Y (nx266), .A0 (nx2580), .A1 (nx2874)) ;
    nor02ii ix209 (.Y (nx208), .A0 (nx2848), .A1 (random_num_input[0])) ;
    nor02ii ix217 (.Y (nx216), .A0 (nx2846), .A1 (random_num_input[1])) ;
    nor02ii ix227 (.Y (nx226), .A0 (nx2840), .A1 (random_num_input[2])) ;
    nor02ii ix235 (.Y (nx234), .A0 (nx2836), .A1 (random_num_input[3])) ;
    nor02ii ix247 (.Y (nx246), .A0 (nx2832), .A1 (random_num_input[4])) ;
    nor02ii ix255 (.Y (nx254), .A0 (nx2830), .A1 (random_num_input[5])) ;
    nor02ii ix345 (.Y (nx344), .A0 (nx2876), .A1 (nx342)) ;
    nor02ii ix277 (.Y (nx276), .A0 (nx2852), .A1 (random_num_input[0])) ;
    nor02ii ix285 (.Y (nx284), .A0 (nx2848), .A1 (random_num_input[1])) ;
    nor02ii ix295 (.Y (nx294), .A0 (nx2846), .A1 (random_num_input[2])) ;
    nor02ii ix303 (.Y (nx302), .A0 (nx2840), .A1 (random_num_input[3])) ;
    nor02ii ix315 (.Y (nx314), .A0 (nx2506), .A1 (random_num_input[6])) ;
    nor02ii ix323 (.Y (nx322), .A0 (nx2836), .A1 (random_num_input[4])) ;
    nor02ii ix331 (.Y (nx330), .A0 (nx2832), .A1 (random_num_input[5])) ;
    nor02ii ix433 (.Y (nx432), .A0 (nx2638), .A1 (nx2874)) ;
    nor02ii ix355 (.Y (nx354), .A0 (nx2856), .A1 (random_num_input[0])) ;
    nor02ii ix363 (.Y (nx362), .A0 (nx2852), .A1 (random_num_input[1])) ;
    nor02ii ix373 (.Y (nx372), .A0 (nx2848), .A1 (random_num_input[2])) ;
    nor02ii ix381 (.Y (nx380), .A0 (nx2846), .A1 (random_num_input[3])) ;
    nor02ii ix393 (.Y (nx392), .A0 (nx2840), .A1 (random_num_input[4])) ;
    nor02ii ix401 (.Y (nx400), .A0 (nx2836), .A1 (random_num_input[5])) ;
    nor02ii ix411 (.Y (nx410), .A0 (nx2515), .A1 (random_num_input[6])) ;
    nor02ii ix419 (.Y (nx418), .A0 (nx2506), .A1 (random_num_input[7])) ;
    nor02ii ix509 (.Y (nx508), .A0 (nx2876), .A1 (nx506)) ;
    nor02ii ix441 (.Y (nx440), .A0 (nx2856), .A1 (random_num_input[1])) ;
    nor02ii ix449 (.Y (nx448), .A0 (nx2852), .A1 (random_num_input[2])) ;
    nor02ii ix459 (.Y (nx458), .A0 (nx2848), .A1 (random_num_input[3])) ;
    nor02ii ix467 (.Y (nx466), .A0 (nx2846), .A1 (random_num_input[4])) ;
    nor02ii ix479 (.Y (nx478), .A0 (nx2515), .A1 (random_num_input[7])) ;
    nor02ii ix487 (.Y (nx486), .A0 (nx2840), .A1 (random_num_input[5])) ;
    nor02ii ix495 (.Y (nx494), .A0 (nx2528), .A1 (random_num_input[6])) ;
    nor02ii ix575 (.Y (nx574), .A0 (nx2700), .A1 (ready_1)) ;
    nor02ii ix517 (.Y (nx516), .A0 (nx2856), .A1 (random_num_input[2])) ;
    nor02ii ix525 (.Y (nx524), .A0 (nx2852), .A1 (random_num_input[3])) ;
    nor02ii ix535 (.Y (nx534), .A0 (nx2848), .A1 (random_num_input[4])) ;
    nor02ii ix543 (.Y (nx542), .A0 (nx2846), .A1 (random_num_input[5])) ;
    nor02ii ix555 (.Y (nx554), .A0 (nx2545), .A1 (random_num_input[6])) ;
    nor02ii ix563 (.Y (nx562), .A0 (nx2528), .A1 (random_num_input[7])) ;
    nor02ii ix631 (.Y (nx630), .A0 (nx2826), .A1 (nx628)) ;
    nor02ii ix583 (.Y (nx582), .A0 (nx2545), .A1 (random_num_input[7])) ;
    nor02ii ix591 (.Y (nx590), .A0 (nx2856), .A1 (random_num_input[3])) ;
    nor02ii ix599 (.Y (nx598), .A0 (nx2852), .A1 (random_num_input[4])) ;
    nor02ii ix609 (.Y (nx608), .A0 (nx2848), .A1 (random_num_input[5])) ;
    nor02ii ix617 (.Y (nx616), .A0 (nx2568), .A1 (random_num_input[6])) ;
    nor02ii ix677 (.Y (nx676), .A0 (nx2743), .A1 (ready_1)) ;
    nor02ii ix639 (.Y (nx638), .A0 (nx2856), .A1 (random_num_input[4])) ;
    nor02ii ix647 (.Y (nx646), .A0 (nx2852), .A1 (random_num_input[5])) ;
    nor02ii ix657 (.Y (nx656), .A0 (nx2588), .A1 (random_num_input[6])) ;
    nor02ii ix667 (.Y (nx666), .A0 (nx2568), .A1 (random_num_input[7])) ;
    nor02ii ix713 (.Y (nx712), .A0 (nx2826), .A1 (nx710)) ;
    nor02ii ix685 (.Y (nx684), .A0 (nx2856), .A1 (random_num_input[5])) ;
    nor02ii ix693 (.Y (nx692), .A0 (nx2615), .A1 (random_num_input[6])) ;
    nor02ii ix703 (.Y (nx702), .A0 (nx2588), .A1 (random_num_input[7])) ;
    nor02ii ix739 (.Y (nx738), .A0 (nx2769), .A1 (ready_1)) ;
    nor02ii ix721 (.Y (nx720), .A0 (nx2646), .A1 (random_num_input[6])) ;
    nor02ii ix729 (.Y (nx728), .A0 (nx2615), .A1 (random_num_input[7])) ;
    nor02ii ix755 (.Y (nx754), .A0 (nx2826), .A1 (row_7_14)) ;
    nor02ii ix747 (.Y (nx746), .A0 (nx2646), .A1 (random_num_input[7])) ;
    or02 ix2813 (.Y (nx2814), .A0 (reset_rows), .A1 (ready_1)) ;
    or02 ix2815 (.Y (nx2816), .A0 (reset_rows), .A1 (ready_1)) ;
    latchs_ni lat_complete_fsm_u1 (.QB (nx5), .D (nx2453), .CLK (nx2860), .S (
              nx2810)) ;
    inv02 lat_complete_fsm_u2 (.Y (complete), .A (nx5)) ;
    latchs_ni lat_reset_rows_u1 (.QB (nx2870), .D (nx2453), .CLK (complete), .S (
              clk)) ;
    inv02 lat_reset_rows_u2 (.Y (reset_rows), .A (nx2870)) ;
    latchs_ni lat_ready_1_u1 (.QB (nx2872), .D (nx2453), .CLK (nx2860), .S (
              nx2860)) ;
    inv02 lat_ready_1_u2 (.Y (ready_1), .A (nx2872)) ;
    inv02 lat_ready_1_u2_rep_1 (.Y (nx2874), .A (nx2872)) ;
    inv01 ix2875 (.Y (nx2876), .A (nx2874)) ;
endmodule

